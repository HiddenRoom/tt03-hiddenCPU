module alu
(
  input [1:0] opcode,
  input [7:0] dIn0,
  input [7:0] dIn1,

  output [7:0] dOut,
  output [7:0] pcInc,
  output carry,
  output borrow
);

endmodule
